`default_nettype none

module unified_buffer(
    input wire clk,
    input wire nrst,
    
    
);

endmodule

`default_nettype wire