`default_nettype none

module TPU(
    input wire clk,
    input wire nrst, 

    // spi interface
);

endmodule

`default_nettype wire