`default_nettype none

module mux #(
    parameter SEL_WIDTH = 1,
    parameter OUT_NUM = 2 ** (SEL_WIDTH)
)(
    
);

endmodule

`default_nettype wire